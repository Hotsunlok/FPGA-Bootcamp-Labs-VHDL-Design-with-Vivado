library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package math_package is
    function AC_COUNTDOWN(curr_value : integer) return integer;
    function FN_COUNTDOWN(curr_value : integer) return integer;
end package math_package;
